library verilog;
use verilog.vl_types.all;
entity top_tb is
    generic(
        period          : integer := 20
    );
end top_tb;
