library verilog;
use verilog.vl_types.all;
entity FSM_Execution_Unit is
    generic(
        G30_1           : integer := 0;
        G30_3           : integer := 1;
        G30_4           : integer := 2;
        G30_5           : integer := 3;
        G30_e           : integer := 4;
        G30_2           : integer := 5;
        RES             : integer := 6;
        G28_1           : integer := 7;
        G28_2           : integer := 8;
        G28_3           : integer := 9;
        G28_5           : integer := 10;
        G28_4           : integer := 11;
        G28_e           : integer := 12;
        G29_1           : integer := 13;
        G29_2           : integer := 14;
        G29_3           : integer := 15;
        G29_5           : integer := 16;
        G29_4           : integer := 17;
        G29_e           : integer := 18;
        FETCH           : integer := 19;
        G1_1            : integer := 20;
        G2_1            : integer := 21;
        G3_1            : integer := 22;
        G4_1            : integer := 23;
        G9_1            : integer := 24;
        G5_1            : integer := 25;
        G6_1            : integer := 26;
        G7_1            : integer := 27;
        G8_1            : integer := 28;
        G19_1           : integer := 29;
        G15_1           : integer := 30;
        G15_3           : integer := 31;
        G15_4           : integer := 32;
        G15_5           : integer := 33;
        G15_2           : integer := 34;
        G15_7           : integer := 35;
        G15_e3          : integer := 36;
        G15_6           : integer := 37;
        G15_e2          : integer := 38;
        G15_e1          : integer := 39;
        G15_8           : integer := 40;
        G10_1           : integer := 41;
        G10_3           : integer := 42;
        G10_4           : integer := 43;
        G10_5           : integer := 44;
        G10_2           : integer := 45;
        G10_7           : integer := 46;
        G10_e3          : integer := 47;
        G10_e1          : integer := 48;
        G10_e2          : integer := 49;
        G10_6           : integer := 50;
        G10_8           : integer := 51;
        G17_1           : integer := 52;
        G17_4           : integer := 53;
        G17_6           : integer := 54;
        G17_3           : integer := 55;
        G17_2           : integer := 56;
        G17_8           : integer := 57;
        G17_9           : integer := 58;
        G17_7           : integer := 59;
        G17_5           : integer := 60;
        G17_10          : integer := 61;
        G17_e           : integer := 62;
        G17_11          : integer := 63;
        G16_1           : integer := 64;
        G16_3           : integer := 65;
        G16_4           : integer := 66;
        G16_5           : integer := 67;
        G16_2           : integer := 68;
        G16_7           : integer := 69;
        G16_6           : integer := 70;
        G16_e3          : integer := 71;
        G16_e1          : integer := 72;
        G16_e2          : integer := 73;
        G16_8           : integer := 74;
        G11_1           : integer := 75;
        G11_5           : integer := 76;
        G11_6           : integer := 77;
        G11_2           : integer := 78;
        G11_7           : integer := 79;
        G11_3           : integer := 80;
        G11_4           : integer := 81;
        G11_e           : integer := 82;
        G31_1           : integer := 83;
        G34_1           : integer := 84;
        G32_1           : integer := 85;
        G33_1           : integer := 86;
        G12_1           : integer := 87;
        G12_e1          : integer := 88;
        G12_e2          : integer := 89;
        G12_2           : integer := 90;
        G12_3           : integer := 91;
        G12_4           : integer := 92;
        G20_1           : integer := 93;
        G20_2           : integer := 94;
        G20_5           : integer := 95;
        G20_e           : integer := 96;
        G20_3           : integer := 97;
        G20_4           : integer := 98;
        G21_1           : integer := 99;
        G21_2           : integer := 100;
        G21_3           : integer := 101;
        G21_4           : integer := 102;
        G21_e           : integer := 103;
        G13_3           : integer := 104;
        G13_1           : integer := 105;
        G13_4           : integer := 106;
        G13_2           : integer := 107;
        G13_e1          : integer := 108;
        G13_e2          : integer := 109;
        G18_1           : integer := 110;
        G18_2           : integer := 111;
        G18_3           : integer := 112;
        G18_4           : integer := 113;
        G18_e           : integer := 114;
        G18_5           : integer := 115;
        G26_1           : integer := 116;
        G26_2           : integer := 117;
        G26_3           : integer := 118;
        G26_4           : integer := 119;
        G26_e           : integer := 120;
        G27_1           : integer := 121;
        G27_2           : integer := 122;
        G27_3           : integer := 123;
        G27_4           : integer := 124;
        G27_e           : integer := 125;
        G14_1           : integer := 126;
        G14_5           : integer := 127;
        G14_6           : integer := 128;
        G14_2           : integer := 129;
        G14_7           : integer := 130;
        G14_3           : integer := 131;
        G14_4           : integer := 132;
        G14_e           : integer := 133;
        G22_1           : integer := 134;
        G22_e           : integer := 135;
        G23_1           : integer := 136;
        G23_e           : integer := 137;
        G24_1           : integer := 138;
        G24_2           : integer := 139;
        G24_e           : integer := 140;
        G25_1           : integer := 141;
        G25_2           : integer := 142;
        G25_e           : integer := 143
    );
    port(
        adr_nxt_pc_i    : in     vl_logic_vector(15 downto 0);
        adr_pc_i        : in     vl_logic_vector(15 downto 0);
        adr_sp_i        : in     vl_logic_vector(15 downto 0);
        alu_dec_val_i   : in     vl_logic_vector(7 downto 0);
        clk_clk_i       : in     vl_logic;
        d_alu_i         : in     vl_logic_vector(7 downto 0);
        d_i             : in     vl_logic_vector(7 downto 0);
        d_regs_out_i    : in     vl_logic_vector(7 downto 0);
        irq_n_i         : in     vl_logic;
        nmi_i           : in     vl_logic;
        q_a_i           : in     vl_logic_vector(7 downto 0);
        q_x_i           : in     vl_logic_vector(7 downto 0);
        q_y_i           : in     vl_logic_vector(7 downto 0);
        rdy_i           : in     vl_logic;
        reg_0flag_i     : in     vl_logic;
        reg_1flag_i     : in     vl_logic;
        reg_7flag_i     : in     vl_logic;
        rst_rst_n_i     : in     vl_logic;
        so_n_i          : in     vl_logic;
        a_o             : out    vl_logic_vector(15 downto 0);
        adr_o           : out    vl_logic_vector(15 downto 0);
        ch_a_o          : out    vl_logic_vector(7 downto 0);
        ch_b_o          : out    vl_logic_vector(7 downto 0);
        d_o             : out    vl_logic_vector(7 downto 0);
        d_regs_in_o     : out    vl_logic_vector(7 downto 0);
        fetch_o         : out    vl_logic;
        ld_o            : out    vl_logic_vector(1 downto 0);
        ld_pc_o         : out    vl_logic;
        ld_sp_o         : out    vl_logic;
        load_regs_o     : out    vl_logic;
        offset_o        : out    vl_logic_vector(15 downto 0);
        rd_o            : out    vl_logic;
        sel_pc_in_o     : out    vl_logic;
        sel_pc_val_o    : out    vl_logic_vector(1 downto 0);
        sel_rb_in_o     : out    vl_logic_vector(1 downto 0);
        sel_rb_out_o    : out    vl_logic_vector(1 downto 0);
        sel_reg_o       : out    vl_logic_vector(1 downto 0);
        sel_sp_as_o     : out    vl_logic;
        sel_sp_in_o     : out    vl_logic;
        sync_o          : out    vl_logic;
        wr_o            : out    vl_logic
    );
end FSM_Execution_Unit;
